package shared_package;
    bit test_finished;
    integer error_count, correct_count;
endpackage